`define KEY = 256'h34d20ac43f554f1d2fd101496787e3954e39d417e33528f13c005501aa1a9e47;
`define IV = 64'hb97b7f467edaefd8;
