`define GOWIN