`define GOWIN
`define INV_PORTS